// Ori in included in the or operation in alu, but multiply is not completed by now.
module cpu (
    input  wire        clk,
    input  wire        resetn,
    // inst sram interface
    output wire        inst_sram_en,
    output wire [31:0] inst_sram_addr,
    input  wire [31:0] inst_sram_rdata,
    // data sram interface
    output wire        data_sram_en,
    output wire [3:0]  data_sram_wen,
    output wire [31:0] data_sram_addr,
    output wire [31:0] data_sram_wdata,
    input  wire [31:0] data_sram_rdata,
    // trace debug interface
    output wire [31:0] debug_wb_pc,
    output wire  debug_wb_rf_wen,
    output wire [ 4:0] debug_wb_rf_wnum,
    output wire [31:0] debug_wb_rf_wdata
);
// signal valid define(use reset instead of resetn)
  reg reset;
  always @(posedge clk) reset <= ~resetn;

  reg valid;
  always @(posedge clk) begin
    if (reset) begin
      valid <= 1'b0;
    end else begin
      valid <= 1'b1;
    end
  end
  assign inst_sram_en = valid;
// signal define
  wire [31:0] seq_pc;
  wire [31:0] nextpc;
  wire        br_taken; // branch taken signal
  wire [31:0] br_target; // branch target address
  wire [31:0] inst; // instruction
  reg  [31:0] pc; // program counter

  wire [11:0] alu_op;
  wire        load_op;
  wire        src2_is_imm; // src2 is immediate number
  wire        res_from_mem; //load is 1, or from alu_result
  wire        gr_we; // no st/b/beq
  wire        mem_we; //store is 1
  wire        src_reg_is_rd; //beq use rd
  wire [ 4:0] dest; // write register address
  wire [31:0] rj_value;
  wire [31:0] rkd_value;
  wire [31:0] imm; // immediate number (extend)
  wire [31:0] br_offs;
// Instruction decode
  wire [ 5:0] op_31_26;
  wire [ 3:0] op_25_22;
  wire [ 1:0] op_21_20;
  wire [ 4:0] op_19_15;
  wire [ 4:0] rd;
  wire [ 4:0] rj;
  wire [ 4:0] rk;
// for instant number
  wire [11:0] i12;
  wire [15:0] i16;
  wire [25:0] i26;
// for decoders.v
  wire [63:0] op_31_26_d;
  wire [15:0] op_25_22_d;
  wire [ 3:0] op_21_20_d;
  wire [31:0] op_19_15_d;

  wire        inst_mul_w;
  wire        inst_add_w;
  wire        inst_sub_w;
  wire        inst_slti;
  wire        inst_and;
  wire        inst_slli_w;
  wire        inst_addi_w;
  wire        inst_ld_w;
  wire        inst_st_w;
  wire        inst_b;
  wire        inst_beq;
  wire        inst_ori;

  wire        need_ui5;
  wire        need_si12;
  wire        need_si16;
  wire        need_si26;
  wire        need_ui12;

  wire [ 4:0] rf_raddr1;
  wire [31:0] rf_rdata1;
  wire [ 4:0] rf_raddr2;
  wire [31:0] rf_rdata2;
  wire        rf_we;
  wire [ 4:0] rf_waddr;
  wire [31:0] rf_wdata;

  wire [31:0] alu_src1;
  wire [31:0] alu_src2;
  wire [31:0] alu_result;
  wire [31:0] mult_result;
  wire [31:0] mem_result;

// PC update (if branch jumping then use br_target, otherwise use seq_pc)
  assign seq_pc = pc + 3'h4;
  assign nextpc = br_taken ? br_target : seq_pc;

  always @(posedge clk) begin
    if (reset) begin
      pc <= 32'hfffffffc;  //trick: to make nextpc be 0x00000000 during reset
    end else begin
      pc <= nextpc;
    end
  end


  assign inst_sram_addr  = pc;
  assign inst            = inst_sram_rdata;

  assign op_31_26        = inst[31:26];
  assign op_25_22        = inst[25:22];
  assign op_21_20        = inst[21:20];
  assign op_19_15        = inst[19:15];

  assign rd              = inst[4:0];
  assign rj              = inst[9:5];
  assign rk              = inst[14:10];

  assign i12             = inst[21:10];
  assign i16             = inst[25:10];
  assign i26             = {inst[9:0], inst[25:10]};

  decoder_6_64 u_dec0 (
      .in (op_31_26),
      .out(op_31_26_d)
  );
  decoder_4_16 u_dec1 (
      .in (op_25_22),
      .out(op_25_22_d)
  );
  decoder_2_4 u_dec2 (
      .in (op_21_20),
      .out(op_21_20_d)
  );
  decoder_5_32 u_dec3 (
      .in (op_19_15),
      .out(op_19_15_d)
  );

  assign inst_add_w = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h00];
  assign inst_sub_w = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h02];
  assign inst_slti = op_31_26_d[6'h00] & op_25_22_d[4'h8];
  assign inst_and = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h09];
  assign inst_slli_w = op_31_26_d[6'h00] & op_25_22_d[4'h1] & op_21_20_d[2'h0] & op_19_15_d[5'h01];
  assign inst_addi_w = op_31_26_d[6'h00] & op_25_22_d[4'ha];
  assign inst_ld_w = op_31_26_d[6'h0a] & op_25_22_d[4'h2];
  assign inst_st_w = op_31_26_d[6'h0a] & op_25_22_d[4'h6];
  assign inst_b = op_31_26_d[6'h14];
  assign inst_beq = op_31_26_d[6'h16];
  assign inst_ori = op_31_26_d[6'h00] & op_25_22_d[4'he];
  // This step is not completed, a multiplier generated by ip core is needed
  assign inst_mul_w = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h18];

  assign alu_op[0] = inst_add_w | inst_addi_w | inst_ld_w | inst_st_w; // add
  assign alu_op[1] = inst_sub_w;  // sub
  assign alu_op[2] = inst_slti;  // slti(need to rewrite)
  assign alu_op[3] = 1'b0;  // ult
  assign alu_op[4] = inst_and;  // and
  assign alu_op[5] = 1'b0;  // nor
  assign alu_op[6] = inst_ori;  // ori(need to rewrite)
  assign alu_op[7] = 1'b0;  // xor
  assign alu_op[8] = inst_slli_w;  // sll
  assign alu_op[9] = 1'b0;  // srl
  assign alu_op[10] = 1'b0;  // sra
  assign alu_op[11] = 1'b0;

  assign need_ui5 = inst_slli_w;
  assign need_ui12 = inst_ori;
  assign need_si12 = inst_addi_w | inst_ld_w | inst_st_w | inst_slti;
  assign need_si16 = inst_beq ;
  assign need_si26 = inst_b ;
//this Line should be rewritten
  assign imm = need_ui5  ? {27'h0, rk[4:0]} :
               need_si12 ? {{20{i12[11]}}, i12[11:0]} :
               need_ui12 ? {20'h0, i12[11:0]} :
               32'h0;

  assign br_offs = need_si26 ? {{4{i26[25]}}, i26[25:0], 2'b0} : {{14{i16[15]}}, i16[15:0], 2'b0};

  assign src_reg_is_rd = inst_beq | inst_st_w;

  assign src2_is_imm   = inst_slli_w |
                       inst_addi_w |
                       inst_ld_w   |
                       inst_st_w   |
                       inst_ori    |
                       inst_slti;

  assign res_from_mem = inst_ld_w;
  assign gr_we = ~inst_st_w & ~inst_beq & ~inst_b;  // ! error
  assign mem_we = inst_st_w;
  assign dest = rd;

  assign rf_raddr1 = rj;
  assign rf_raddr2 = src_reg_is_rd ? rd : rk;
  reg_file u_regfile (
      .clk   (clk),
      .raddr1(rf_raddr1),
      .rdata1(rf_rdata1),
      .raddr2(rf_raddr2),
      .rdata2(rf_rdata2),
      .we    (rf_we),
      .waddr (rf_waddr),
      .wdata (rf_wdata)
  );

  assign rj_value  = rf_rdata1;
  assign rkd_value = rf_rdata2;

  wire rj_eq_rd = (rj_value == rkd_value);  // ! error
  assign br_taken = (   inst_beq  &&  rj_eq_rd
                   || inst_b
                  ) && valid;
  assign br_target = pc + br_offs; 

  assign alu_src1 =  rj_value;
  assign alu_src2 = src2_is_imm ? imm : rkd_value;

  simple_alu u_alu (
      .alu_op    (alu_op),
      .alu_src1  (alu_src1),   // ! error
      .alu_src2  (alu_src2),
      .alu_result(alu_result)
  );
  multi u_multi (
      .multiplicand(alu_src1),
      .multiplier(alu_src2),
      .product_low(mult_result)
  );
  assign data_sram_en =  (inst_st_w | inst_ld_w) && valid;
  assign data_sram_wen = (mem_we && valid) ? 4'b1111 : 4'b0000;
  assign data_sram_addr  = (inst_st_w | inst_ld_w) ? alu_result : 32'b0; // ! warn: addr out of bound
  assign data_sram_wdata = rkd_value;

  assign mem_result = data_sram_rdata;
  wire [31:0] final_result = res_from_mem ? mem_result : inst_mul_w ? mult_result : alu_result;  // ! error

  assign rf_we             = gr_we && valid && (dest != 5'b00000);
  assign rf_waddr          = dest;
  assign rf_wdata          = final_result;

  // debug info generate
  assign debug_wb_pc       = pc;
  assign debug_wb_rf_wen   = rf_we;
  assign debug_wb_rf_wnum  = dest;
  assign debug_wb_rf_wdata = final_result;

endmodule