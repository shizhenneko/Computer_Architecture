module id_stage(
    input clk,
    input resetn,
// control signal between id if exe
    output id_allow_in,
    input if_to_id_valid,
    input exe_allow_in,
    output id_to_exe_valid,
// hazard detection
    input exe_rf_we,
    input [4:0] exe_rf_waddr,
    input [31:0] exe_rf_wdata,
    input exe_valid,
    input mem_rf_we,
    input [4:0] mem_rf_waddr,
    input [31:0] mem_rf_wdata,
    input mem_valid,
    input wb_valid,
    input exe_is_load,
// if send to id for pc update
    input [31:0] if_pc,
    input [31:0] inst,
// id sent to if for branch selection
    output br_taken,
    output br_cancel,
    output [31:0] br_target,
// if send to exe
    output [31:0] rj_value,
    output [31:0] rkd_value,
    output [31:0] imm,
    output [11:0] alu_op,
    output src2_is_imm,
    output res_from_mem,
    output reg_we,
    output id_is_multi,
    output mem_en,
    output [3:0] mem_we,
    output [4:0] reg_waddr,
// wb send to id  for regfile
    input wb_rf_we,
    input [4:0] wb_rf_waddr,
    input [31:0] wb_rf_wdata,
// expose latched pc to next stage
    output [31:0] id_pc
);
    wire reset = ~resetn;
// pipeline register
    reg [31:0] id_pc;
    reg [31:0] id_inst;
// input bus from wb
    // use inputs directly: wb_rf_we, wb_rf_waddr, wb_rf_wdata

// output to exe
    // driven via assigns to output ports
// output to if
    // use output ports directly: br_taken, br_cancel
//control signal
    reg id_valid;
    wire id_ready_go;

// signal assignment
    assign id_allow_in = !id_valid || (id_ready_go && exe_allow_in);
    assign id_to_exe_valid = id_valid && id_ready_go;
// pipeline update logic
    always @(posedge clk) begin
        if (reset) begin
            id_valid <= 1'b0;
        end else if (br_cancel) begin
            id_valid <= 1'b0;
        end else if (id_allow_in) begin
            id_valid <= if_to_id_valid;
        end
    end

    always @(posedge clk) begin
        if (id_allow_in && if_to_id_valid) begin
            id_pc <= if_pc;
            id_inst <= inst;
        end
    end
// bypass signal
    // use input exe_rf_waddr directly

// The last thing need to do is to finish the decode
    wire src_reg_is_rd;
    
    wire [5:0] op_31_26;
    wire [3:0] op_25_22;
    wire [1:0] op_21_20;
    wire [4:0] op_19_15;

    wire [4:0] rd;
    wire [4:0] rj;
    wire [4:0] rk;

    wire [11:0] i12;
    wire [15:0] i16;
    wire [25:0] i26;

    wire inst_add_w;
    wire inst_mul_w;
    wire inst_sub_w;
    wire inst_slti;
    wire inst_and;
    wire inst_slli_w;
    wire inst_addi_w;
    wire inst_ld_w;
    wire inst_st_w;
    wire inst_b;
    wire inst_beq;
    wire inst_ori;

    wire need_ui5;
    wire need_si12;
    wire need_si16;
    wire need_si26;
    wire need_ui12;

    wire [ 4:0] rf_raddr1;
    wire [31:0] rf_rdata1;
    wire [ 4:0] rf_raddr2;
    wire [31:0] rf_rdata2;
    wire        rf_we;
    wire [ 4:0] rf_waddr;
    wire [31:0] rf_wdata;

    wire [63:0] op_31_26_d;
    wire [15:0] op_25_22_d;
    wire [ 3:0] op_21_20_d;
    wire [31:0] op_19_15_d;

    assign op_31_26        = inst[31:26];
    assign op_25_22        = inst[25:22];
    assign op_21_20        = inst[21:20];
    assign op_19_15        = inst[19:15];

    assign rd              = inst[4:0];
    assign rj              = inst[9:5];
    assign rk              = inst[14:10];

    assign i12             = inst[21:10];
    assign i16             = inst[25:10];
    assign i26             = inst[25:0];

    decoder_6_64 u_dec0 (
        .in (op_31_26),
        .out(op_31_26_d)
    );
    decoder_4_16 u_dec1 (
        .in (op_25_22),
        .out(op_25_22_d)
    );
    decoder_2_4 u_dec2 (
        .in (op_21_20),
        .out(op_21_20_d)
    );
    decoder_5_32 u_dec3 (
        .in (op_19_15),
        .out(op_19_15_d)
    );

    assign inst_add_w = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h00];
    assign inst_sub_w = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h02];
    assign inst_slti = op_31_26_d[6'h00] & op_25_22_d[4'h8];
    assign inst_and = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h09];
    assign inst_slli_w = op_31_26_d[6'h00] & op_25_22_d[4'h1] & op_21_20_d[2'h0] & op_19_15_d[5'h01];
    assign inst_addi_w = op_31_26_d[6'h00] & op_25_22_d[4'ha];
    assign inst_ld_w = op_31_26_d[6'h0a] & op_25_22_d[4'h2];
    assign inst_st_w = op_31_26_d[6'h0a] & op_25_22_d[4'h6];
    assign inst_b = op_31_26_d[6'h14];
    assign inst_beq = op_31_26_d[6'h16];
    assign inst_ori = op_31_26_d[6'h00] & op_25_22_d[4'he];
    // This step is not completed, a multiplier generated by ip core is needed
    assign inst_mul_w = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h18];

    assign alu_op[0] = inst_add_w | inst_addi_w | inst_ld_w | inst_st_w; // add
    assign alu_op[1] = inst_sub_w;  // sub
    assign alu_op[2] = inst_slti;  // slti(need to rewrite)
    assign alu_op[3] = 1'b0;  // ult
    assign alu_op[4] = inst_and;  // and
    assign alu_op[5] = 1'b0;  // nor
    assign alu_op[6] = inst_ori;  // ori(need to rewrite)
    assign alu_op[7] = 1'b0;  // xor
    assign alu_op[8] = inst_slli_w;  // sll
    assign alu_op[9] = 1'b0;  // srl
    assign alu_op[10] = 1'b0;  // sra
    assign alu_op[11] = 1'b0;

    assign need_ui5 = inst_slli_w;
    assign need_ui12 = inst_ori;
    assign need_si12 = inst_addi_w | inst_ld_w | inst_st_w | inst_slti;
    assign need_si16 = inst_beq ;
    assign need_si26 = inst_b ;
    //this Line should be rewritten
    assign imm = need_ui5  ? {27'h0, rk[4:0]} :
                need_si12 ? {{20{i12[11]}}, i12[11:0]} :
                need_ui12 ? {20'h0, i12[11:0]} :
                32'h0;

    wire [31:0] br_offs;
    assign br_offs = need_si26 ? {{4{i26[25]}}, i26[25:0], 2'b0} : {{14{i16[15]}}, i16[15:0], 2'b0};

    assign src_reg_is_rd = inst_beq | inst_st_w;
    assign br_target = id_pc + br_offs;

    assign src2_is_imm   = inst_slli_w |
                        inst_addi_w |
                        inst_ld_w   |
                        inst_st_w   |
                        inst_ori    |
                        inst_slti;
    assign res_from_mem = inst_ld_w;
    assign reg_we = id_valid & (rd != 5'd0) & ~inst_st_w & ~inst_beq & ~inst_b;
    assign mem_en = inst_ld_w | inst_st_w;
    assign mem_we = {4{inst_st_w}};
    assign reg_waddr = rd;
    assign id_is_multi = inst_mul_w;
    assign rf_raddr1 = rj;
    assign rf_raddr2 = src_reg_is_rd ? rd : rk;    

reg_file u_reg_file (
    .clk (clk),
    .raddr1 (rf_raddr1),
    .raddr2 (rf_raddr2),
    .waddr (rf_waddr),
    .wdata (rf_wdata),
    .we (rf_we),
    .rdata1 (rf_rdata1),
    .rdata2 (rf_rdata2)
);
    // forwarding will drive rj_value and rkd_value below

    wire rj_eq_rd = (rj_value == rkd_value);
    assign br_taken = id_valid && ( inst_beq && rj_eq_rd || inst_b) && id_ready_go;
// pass hazard from wb
    assign rf_we = wb_rf_we;
    assign rf_waddr = wb_rf_waddr;
    assign rf_wdata = wb_rf_wdata;
// when RAW may happen
    wire use_rf_rdata1 = id_valid && !inst_b;
    wire use_rf_rdata2 = id_valid && (inst_add_w || inst_sub_w || inst_slti || inst_and || inst_beq || inst_mul_w || inst_st_w);
// hazard
wire rf_rdata1_hazard = use_rf_rdata1 && (exe_valid && exe_is_load && exe_rf_we && (rf_raddr1 == exe_rf_waddr));
wire rf_rdata2_hazard = use_rf_rdata2 && (exe_valid && exe_is_load && exe_rf_we && (rf_raddr2 == exe_rf_waddr));
assign id_ready_go = !rf_rdata1_hazard && !rf_rdata2_hazard;

assign br_cancel = id_valid && br_taken && id_ready_go && exe_allow_in;

assign rj_value = (exe_valid && exe_rf_we && (rf_raddr1 == exe_rf_waddr)) ? exe_rf_wdata : (mem_valid && mem_rf_we && (rf_raddr1 == mem_rf_waddr)) ? mem_rf_wdata : (wb_valid && wb_rf_we && (rf_raddr1 == wb_rf_waddr)) ? wb_rf_wdata : rf_rdata1;

assign rkd_value = (exe_valid && exe_rf_we && (rf_raddr2 == exe_rf_waddr)) ? exe_rf_wdata : (mem_valid && mem_rf_we && (rf_raddr2 == mem_rf_waddr)) ? mem_rf_wdata : (wb_valid && wb_rf_we && (rf_raddr2 == wb_rf_waddr)) ? wb_rf_wdata : rf_rdata2;

endmodule